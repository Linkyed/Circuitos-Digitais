module decisor (A, B, out);

   input   A, B; // ENTRADAS DO MODULO RELACIONADA A ATIVAÇÃO DA FUNÇÃO DOIS EM CADA DAS INTERFACES
   output  [1:0] out; // SAIDAS DO MODULO RELACIONADAS A SE A FUNCIONALIDADE 2 FOI ATIVADA, E QUAL DAS DUAS INTERFACES
							 // DEVE TER SEU CODIGO PASSADO (1 PARA A IE02 TER SEU CODIGO PASSADO E 0 PARA A IE01 TER SEU CODIGO PASSADO PARA FRENTE)
	 
	// PORTAS LOGICAS OR PARA GERAR AS DUAS SAIDAS DO MODULO
	or out0 (out[0], A, B);
	or out1 (out[1], A);

endmodule