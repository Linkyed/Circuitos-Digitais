module FUN2_P_S(A, B, C, D, E, F, out);
   input A, B, C, D, E, F;
   output [2:0] out;
	
	xor Xor0 (out[0], A, D);
	xor Xor1 (out[1], B, E);
	xor Xor2 (out[2], C, F);

	
endmodule