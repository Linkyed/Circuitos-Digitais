module conv_per_bin(A, B, C, out);
   input A, B, C; // ENTRADAS DO MODULO RELACIONADA AS CHAVES QUE DETERMINAM O PERFIL DA INTERFACE
   output [1:0] out; // SAIDA DO MODULO RELACIONADA AO BINARIO DE 2 BITS GERADO ATRAVES DO CODIGO DO PERFIL
	
	wire A_not, B_not,// FIO PARA SER UTILIZADO EM UM PORTA INVERSORA
	SUP1, SUP2; // FIOS DE SUPORTE PARA SEREM USADOS EM PORTAS LOGICAS
	
	//PORTAS INVERSORAS PARA AS ENTRADAS A e B
	not A_inv (A_not, A);
	not B_inv (B_not, B);
	
	//PORTAS LOGICAS INTERMEDIARAS PARA TEREM SUAS SAIDAS UTILIZADAS NO OUTPUT DO MODULO
	and And3 (SUP1, A_not, B, C);
	and And2 (SUP2, A, B_not, C); 
	
	//SAIDAS QUE REPRESENTARÃO O PERFIL EM BINARIO DE 2 DIGITOS SEGUINDO A ORDEM:
   //(ADM = 11, TESTER = 10, USER = 01, GUEST = 00)
	or Or0 (out[0], SUP1, SUP2);
	and And0 (out[1], C, B_not);
	
endmodule