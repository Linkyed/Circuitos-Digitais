module TESTES( LED0, LED2, LED3, LED5, 
					M_LED0, M_LED1, M_LED2, M_LED3, M_LED4, M_LED5, M_LED6, MCOL_LED0,
					RGB_r,
					CH7, CH6, CH5, CH4, B3, B2, 
					CH3, CH2, CH1, CH0, B1, B0, 
					SEG7_a, SEG7_b, SEG7_c, SEG7_d, SEG7_e, SEG7_f, SEG7_g, SEG_DP,DITOGO_1,DITIGO_2,DITIGO_3); 
					
   input CH7, CH6, CH5, CH4, B3, B2, // INPUTS DA INTERFACE DE ENTRADA IE01
			CH3, CH2, CH1, CH0, B1, B0; // INPUTS DA INTERFACE DE ENTRADA IE02
			
   output LED0, LED2, LED3, LED5, // OUTPUTS DA INTERFACE DE SAIDA IS02
			 RGB_r, // OUTPUT PARA O LED RGB (VERMELHO)
			 M_LED0, M_LED1, M_LED2, M_LED3, M_LED4, M_LED5, M_LED6, MCOL_LED0, // OUTPUTS DA INTERFACE DE SAIDA IS01
			 SEG7_a, SEG7_b, SEG7_c, SEG7_d, SEG7_e, SEG7_f, SEG7_g,SEG_DP,DITOGO_1,DITIGO_2,DITIGO_3; // OUTPUTS DA INTERFACE DE SAIDA IS03
	
	// FIOS DE 2 BITS PARA:
	wire [1:0] BIN_IE01, BIN_IE02, // CONVERSÃO DO PERFIL EM BINARIO
	SEG7_atv_per; //
	// FIOS DE 3 BITS PARA:
	wire [2: 0] FUN_IE01, FUN_IE02, // ENCAMINHAR A FUNCIONALIDADE ESCOLHIDA PELA INTERFACE
	LEDs_IE01, MATRIZ_IE01, LEDs_IE02, MATRIZ_IE02; // ENCAMINHAR A FUNCIONALIDADE PARA OS DECODIFICADORES
	// FIOS DE 1 BIT PARA: 
	wire PRIO, PRIO_not, // ENCAMINHAR A PRIORIDADE EM RELAÇÃO AOS PERFIS ATUAIS 
	FUN_IGUAIS, // ENCAMINHAR A IGUALDADE ENTRE AS FUNCIONALIDADES SELECIONADAS
	atv_PRIO_IE01, atv_PRIO_IE02, // ENCAMINHAR A ATIVAÇÃO NO CASO DELA SER NECESSARIA
	SEG7_IE01, SEG7_IE02, // ENCAMINHAR A ESCOLHA DA FUNCIONALIDADE 2 PELA INTERFACE
	P_SEG7_0, P_SEG7_1, P_SEG7_2, // ENCAMINHAR O CODIGO DO PERFIL PARA O DECODIFICADOR DE 7 SEGMENTOS
	ver_PIE01, ver_PIE02; // ENCAMINHAR A VERIFICAÇÃO DO PERFIL PARA ACENDER O LED DO PILOTO AUTOMATICO

	// MODULOS RESPONSAVEIS PELA CONVERSÃO DO PERFIL EM BINARIO DE 2 DIGITOS
	conv_per_bin conv_IE01 (CH7, CH6, CH5, BIN_IE01);
	conv_per_bin conv_IE02 (CH3, CH2, CH1, BIN_IE02);
	
	// MODULOS RESPONSAVEIS PELA VALIDAÇÃO DA FUNCIONALIDADE ESCOLHIDA COM BASE NO NIVEL DE ACESSO DO PERFIL ESCOLHIDO
	ver_fun ver_funIE01(FUN_IE01, CH7, CH6, CH5, CH4, B3, B2);
	ver_fun ver_funIE02(FUN_IE02, CH3, CH2, CH1, CH0, B1, B0);
	
	// MODULO PARA COMPARAR AS FUNÇÕES E PERCEBER SE ELAS SÃO IGUAIS OU NÃO
	comp_FUN comp_FUN (FUN_IE01[0], FUN_IE01[1], FUN_IE01[2], FUN_IE02[0], FUN_IE02[1], FUN_IE02[2], FUN_IGUAIS);
	
	// MODULO PARA COMPARAR OS BINARIOS E DECIDIR QUAL DOS DOIS TEM MAIOR PRIORIDADE
	comp_prio comp_prio (BIN_IE01, BIN_IE02, PRIO); 
	
	// PORTA INVERSORA PARA INVERTER A PRIORIDADE PARA IE02 JÁ QUE A PRIORIDADE FUNCIONA DE FORMA INVERÇA PARA ESSA INTERFACE
	not inv_PRIO (PRIO_not, PRIO);
	
	// MODULOS PARA DECIDIR A ATIVAÇÃO DA PRIORIDADE ENTRE AS INTERFACES
	atv_PRIO atv_PRIO0 (PRIO, FUN_IGUAIS, atv_PRIO_IE01);
	atv_PRIO atv_PRIO1 (PRIO_not, FUN_IGUAIS, atv_PRIO_IE02);

	// MODULOS PARA ENCAMINHAR AS FUNCIONALIDADES PARA SEUS DEVIDOS DECODIFICADORES, E TAMBEM RECONHECER A ATIVAÇÃO
	// DA PRIORIDADE
	enc_FUN enc_IE01 (FUN_IE01[0], FUN_IE01[1], FUN_IE01[2], atv_PRIO_IE01, BIN_IE01[0], LEDs_IE01, MATRIZ_IE01, SEG7_IE01);
	enc_FUN enc_IE02 (FUN_IE02[0], FUN_IE02[1], FUN_IE02[2], atv_PRIO_IE02, BIN_IE02[0], LEDs_IE02, MATRIZ_IE02, SEG7_IE02);
	
	// MODULO PARA DECIDIR QUAL DAS DUAS INTERFACES TERA SEU PERFIL APRESENTADO NO MOSTRADOR DE 7 SEGMENTOS
	decisor decisor (SEG7_IE01, SEG7_IE02, SEG7_atv_per);
	
	// MODULO PARA ENCAMINHAR O CODIGO DO PERFIL PARA O MOSTRADOR DE 7 SEGMENTOS
	enc_perf enc_p_0 (CH7, CH3, SEG7_atv_per[0], SEG7_atv_per[1], P_SEG7_0);
	enc_perf enc_p_1 (CH6, CH2, SEG7_atv_per[0], SEG7_atv_per[1], P_SEG7_1);
	enc_perf enc_p_2 (CH5, CH1, SEG7_atv_per[0], SEG7_atv_per[1], P_SEG7_2);
	
	// MODULO DECODIFICADOR PARA MANIPULAR OS LEDS
	decod_Leds Ligar_Leds(LEDs_IE01[0], LEDs_IE01[1], LEDs_IE01[2],LEDs_IE02[0], LEDs_IE02[1], LEDs_IE02[2], LED0, LED2, LED3, LED5);
	
	// MODULO DECODIFICADOR PARA MANIPULAR A MATRIZ DE LEDS 
	wire MCOL_LED0 = 1;
	decod_Matriz Ligar_MLeds(MATRIZ_IE01[0], MATRIZ_IE01[1], MATRIZ_IE01[2],MATRIZ_IE02[0], MATRIZ_IE02[1], MATRIZ_IE02[2], M_LED0, M_LED2, M_LED3, M_LED4 , M_LED5, M_LED6);
	
	// MODULO DECODIFICADOR PARA MANIPULAR O MOSTRADOR DE 7 SEGMENTOS
	wire SEG_DP = 1;
	wire M_LED1 = 1;
	wire DITOGO_1 = 1;
	wire DITIGO_2 = 1;
	wire DITIGO_3 = 1;
	decod_7seg Ligar_7seg (SEG7_a, SEG7_b, SEG7_c, SEG7_d, SEG7_e, SEG7_f, SEG7_g, P_SEG7_0, P_SEG7_1, P_SEG7_2);
	
	// MODULOS PARA VERIFICAR A VALIDADE DO PERFIL SELECIONADO NA INTERFACE
	ver_perf verf_p_IE01 (CH7, CH6, CH5, ver_PIE01);
	ver_perf verf_p_IE02 (CH3, CH2, CH1, ver_PIE02);
	
	// PORTA NOR PARA ACENDER O LED NO CASO EM QUE NÃO EXISTE PERFIL VALIDO EM AMBAS AS INTERFACES
	// E ASSIM DEIXANDO CLARO O FUNCIONAMENTO DO PILOTO AUTOMATICO
	nor (RGB_r, ver_PIE01, ver_PIE02);

endmodule