module ver_perf(A, B, C, out);
   input A, B, C; // ENTRADAS DO MODULO PARA RECEBER AS CHAVES RELACIONADAS AO PERFIL
   output out; // SAIDA DO MODULO QUE RESULTA EM 1 CASO O PERFIL SELECIONADO SEJA UM DOS 4 POSSIVEIS (ADM, TESTER, USER, GUEST)
					// E RESULTA EM 0 CASO O EPRFIL SELECIONADO NÃO SEJA VALIDO
	
	wire A_not, B_not, C_not, // FIOS PARA PORTAS INVERSORAS
	SUP1, SUP2, SUP3, SUP4; // FIOS DE SUPORTE PARA SEREM USADOS EM PORTAS LOGICAS
	
	// PORTAS INVERSORAS PARA TODAS AS ENTRADAS
	not A_inv (A_not, A);
	not B_inv (B_not, B);
	not C_inv (C_not, C);
	
	// SEQUENCIA DE PORTAS LOGICAS PARA VERIFICAR A VALIDADE DO PERFIL(ENTRADAS) INSERIDO NO MODULO
	and And0 (SUP1, A, B_not, C);
	and And1 (SUP2, A_not, B, C);
	and And2 (SUP3, A_not, B_not, C);
	and And3 (SUP4, A, B, C_not);
	
	// PORTA LOGICA OR PARA A SAIDA DO MODULO
	or Or0 (out, SUP1, SUP2, SUP3, SUP4);
	

endmodule