module atv_PRIO (PRIO, FUN_IG, out);
   input PRIO, FUN_IG; // ENTRADAS DO MODULO RELACIONADAS A PRIORIDADE ENTRE OS PERFIS E SE AS FUNCIONALIDADES ESCOLHIDAS FORAM IGUAIS
   output out; // SAIDA DO MODULO RELACIONADA A SE A PRIORIDADE VAI SER ATIVADA OU NÃO NO MODULO
	wire FUN_IG_not; // FIO USADO PARA INVERSÃO DO VALOR DA ENTRADA DE FUNCIONALIDADES IGUAIS
	
	// PORTA INVERSORA PARA A ENTRADA FUN_IG
	not FUN_IG_inv (FUN_IG_not, FUN_IG);
	
	// PORTA LOGICA OR PARA GERAR A UNICA SAIDA DO MODULO
	or Out (out, FUN_IG_not, PRIO);
	
endmodule