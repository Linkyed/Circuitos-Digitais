module enc_FUN(A, B, C, atv_PRIO, INTERF, out_LEDS, out_MATRIZ, out_7SEG);
   input A, B, C, atv_PRIO, INTERF; // ENTRADAS DO MODULO RELACIONADAS A FUNCIONALIDADE ESCOLHIDA PELA INTERFACE,
												// SE A PRIORIDADE TA SENDO ATIVADA OU NÃO E EM QUAL INTERFACE DE SAIDA A FUNCIONALIDADE DEVES SER MOSTRADA
												// INTERF = INTERFACE, E SE FOR 0 SIGNIFICA LEDS E SE FOR 1 MATRIZ
	output [2:0] out_LEDS, out_MATRIZ; // SAIDA DO MODULO QUE APENAS COPIAM A ENTRADA CASO A PRIORIDADE NÃO ESTEJA SENDO
												  // UTILIZADA OU A INTERFACE GANHOU A PRIORIDADE
												  // 3 BITS VÃO PARA O DECODIFICADOR DOS LEDS E OS OUTROS 3 BITS VÃO PARA MATRIZ DE LEDS
	output out_7SEG; // SAIDA RELACIONADA A ATIVAÇÃO DA FUNCIONALIDADE 2
	
	wire INTERF_not, A_not, C_not, // FIOS USADOS PELAS PORTAS INVERSORAS COMO SAIDA
	SUP0, SUP1, SUP2; // FIOS DE SUPORTE PARA AS PORTAS LOGICAS INTERMEDIARIAS
	
	
	// PORTAS INVERSORAS PARA AS ENTRADAS DE INTERFACE, A E C
	not INTERF_inv (INTERF_not, INTERF);
	not A_inv (A_not, A);
	not C_inv (C_not, C);
	
	// PORTAS LOGICAS PARA CRIAR A SAIDA DE 3 BITS QUE SERA LIGADA NO DECODIFICADOR DOS LEDS
	and outLED0 (out_LEDS[0], INTERF_not, A, atv_PRIO);
	or Or0 (SUP0, A, C);
	and outLED1 (out_LEDS[1], INTERF_not, B, atv_PRIO, SUP0);
	and outLED2 (out_LEDS[2], INTERF_not, C, atv_PRIO);	
	
	// PORTAS LOGICAS PARA CRIAR A SAIDA DE 3 BITS QUE SERA LIGADA NO DECODIFICADOR DA MATRIZ DE LEDS
	and outMATRIZ0 (out_MATRIZ[0], INTERF, A, atv_PRIO);
	and And0 (SUP1, B, C, INTERF, atv_PRIO);
	and And1 (SUP2, A, B, INTERF, atv_PRIO);
	or outMATRIZ1 (out_MATRIZ[1], SUP1, SUP2);
	and outMATRIZ2 (out_MATRIZ[2], INTERF, C, atv_PRIO);

	// PORTA LOGICA AND PARA GERAR A SAIDA DA ATIVAÇÃO DA FUNCIONALIDADE 2
	and out7SEG (out_7SEG, A_not, B, C_not, atv_PRIO);
	
endmodule