module comp_FUN(A, B, C, D, E, F, out);
   input A, B, C, D, E, F; // ENTRADAS DO MODULO RELACIONADAS A AMBAS FUNCIONALIDADES DE 3 BITS ESCOLHIDAS PELA INTERFACE
   output out; // SAIDA DO MODULO RELACIONADA A SE AS FUNCIONALIDADES SÃO IGUAIS OU NÃO
	wire igual_0, igual_1, igual_2; // FIOS DE SUPORTE PARA SEREM USADOS NAS PORTAS LOGICAS INTERMEDIARIAS
	
	// PORTAS LOGICAS XNOR PARA VERIFICAR A IGULDADE DE CADA BIT DE UM ENTRADA EM RELAÇÃO A OUTRA
	xnor Or0 (igual_0, A, D);
	xnor Or1 (igual_1, B, E);
	xnor Or2 (igual_2, C, F);
	
	
	// PORTA LOGICA AND PARA GERAR A SAIDA SE AS FUNCIONALIDADES SÃO IGUAIS OU NÃO
	and is_IGUAL (out, igual_0, igual_1, igual_2);
	
endmodule