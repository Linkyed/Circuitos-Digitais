//module atv_PRIO (FUN_IG, PRIO, out);
//   input FUN_IG, PRIO;
//   output [1:0] out;
//	
//	wire out[0] = FUN_IG;
//	
//	
//	
//endmodule