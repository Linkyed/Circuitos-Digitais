module enc_perf (A, B, C, D, out);

   input   A, B, C, D; //ENTRADAS DO MODULO RELACIONADAS AOS BITS DE MESMA SIGNIFICANCIA DE AMBAS INTERFACES,
							  // E TAMBEM RELACIONADA A ATIVAÇÃO DA FUNCONALIDADE 2 E A QUAL VALOR DAS CHAVES DEVE PASSAR PARA A SAIDA DO MODULO
   output  out; // SAIDA DO MODULO RELACIONADA AO VALOR DE QUAL CHAVE DEVE SER PASSADO PARA SAIDA OU SEMPRE 0 CASO
					 // A FUNCIONALIDADE 2 NÃO ESTEJA SENDO ATIVADA
	wire D_not, // FIO USADO NA INVERSÃO DA ENTRADA D
	SUP1, SUP2; // FIOS DE SUPORTE USADOS NAS PORTAS LOGICAS INTERMEDIARIAS
 
	// PORTA INVERSORA PARA ENTRADA D
	not D_inv (D_not, D);
	
	// PORTAS LOGICAS INTERMEDIARIAS PARA SEREM USADAS NA PORTA LOGICA QUE GERA O OUTPUT DO MODULO
   or Or0 (SUP1, A, D);
	or	Or1 (SUP2, B, D_not);
	
	// PORTA LOGICA AND UTILIZADA PARA CONCEDER O OUTPUT DO MODULO
	and And0 (out, C, SUP1, SUP2);

endmodule